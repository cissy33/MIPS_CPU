library verilog;
use verilog.vl_types.all;
entity ram_writefirst_tb is
end ram_writefirst_tb;

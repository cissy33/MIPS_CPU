library verilog;
use verilog.vl_types.all;
entity sltsltu_tb is
end sltsltu_tb;

library verilog;
use verilog.vl_types.all;
entity log_tb is
end log_tb;

library verilog;
use verilog.vl_types.all;
entity pipe_if_tb is
end pipe_if_tb;

library verilog;
use verilog.vl_types.all;
entity bshifter32_carry_tb is
end bshifter32_carry_tb;

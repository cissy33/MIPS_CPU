library verilog;
use verilog.vl_types.all;
entity top_mem_tb is
end top_mem_tb;
